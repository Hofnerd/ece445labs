----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 07/05/2018 04:41:00 PM
-- Design Name: 
-- Module Name: mux2x1 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mux2x132bit is
  Port ( d1, d2 : in std_logic_vector(31 downto 0);
         sel : in std_logic;
         dout : out std_logic_vector(31 downto 0));
end mux2x132bit;

architecture Behavioral of mux2x132bit is

begin

with sel select 
    dout <= d1 when '0',
            d2 when '1',
            X"00000000" when others;
            

end Behavioral;
