library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity pc is

end pc;

architecture behavior of pc is

begin

end behavior;