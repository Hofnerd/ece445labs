library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ALUcntl is
    Port ( Fn   : in STD_LOGIC_VECTOR (5 downto 0);
           Cntl : out STD_LOGIC_VECTOR (3 downto 0));
end ALUcntl;

architecture Behavioral of ALUcntl is

begin

    with Fn select Cntl <=
        "0010" when X"20", --add
        "0010" when X"21", --addu
        "0110" when X"22", --sub
        "0110" when X"23", --subu
        "0000" when X"24", --and
        "0001" when X"25", --or
        "0011" when X"26", --xor
        "1100" when X"27", --nor
        "1111" when X"2A", --slt
        "1110" when X"2B", --sltu
        "0000" when others;

end Behavioral;
